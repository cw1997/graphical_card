library verilog;
use verilog.vl_types.all;
entity graphics_card_vlg_vec_tst is
end graphics_card_vlg_vec_tst;
